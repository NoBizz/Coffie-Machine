module inv(input a, output wire y);

assign y = ~a;

endmodule
